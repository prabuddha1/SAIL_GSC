// key= 10100010
module c1355 (keyInPseudo,  keyIn,  G1,  G10,  G11,  G12,  G13,  G14,  G15,  G16,  G17,  G18,  G19,  G2,  G20,  G21,  G22,  G23,  G24,  G25,  G26,  G27,  G28,  G29,  G3,  G30,  G31,  G32,  G33,  G34,  G35,  G36,  G37,  G38,  G39,  G4,  G40,  G41,  G5,  G6,  G7,  G8,  G9,  G1324,  G1325,  G1326,  G1327,  G1328,  G1329,  G1330,  G1331,  G1332,  G1333,  G1334,  G1335,  G1336,  G1337,  G1338,  G1339,  G1340,  G1341,  G1342,  G1343,  G1344,  G1345,  G1346,  G1347,  G1348,  G1349,  G1350,  G1351,  G1352,  G1353,  G1354,  G1355 ); 
input [7:0] keyIn; 
input  [7:0] keyInPseudo; 
input G1, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9; 
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355; 
wire   N388, N395, N396, N397, N404, N405, N406, N407, N409, N413, n17678, n17679, n17680, n17681, n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689, n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697, n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705, n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713, n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721, n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729, n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737, n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745, n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753, n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761, n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769, n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777, n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785, n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793, n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801, n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809, n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817, n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825, n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833, n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841, n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849; 
assign G1335 = N395;
assign G1336 = N396;
assign G1337 = N397;
assign G1344 = N404;
assign G1345 = N405;
assign G1346 = N406;
assign G1353 = N413;
assign G1338 = n17749z_inv_wire;
XOR2X1 U211 ( .A(n195), .B(n196), .Y(n17749z_inv_wire) );
XOR2X1 U212 ( .A(keyIn[2]), .B(G15), .Y(n196) );
NOR2X1 U213 ( .A(n197), .B(n198), .Y(n195) );
XOR2X1 U214 ( .A(n199), .B(n200), .Y(N413) );
NOR2X1 U215 ( .A(n201), .B(n202), .Y(n200) );
XOR2X1 U216 ( .A(n203), .B(n204), .Y(N406) );
NOR2X1 U217 ( .A(n205), .B(n206), .Y(n204) );
XOR2X1 U218 ( .A(n207), .B(n208), .Y(N405) );
NOR2X1 U219 ( .A(n201), .B(n206), .Y(n208) );
XOR2X1 U220 ( .A(n209), .B(n210), .Y(N404) );
NOR2X1 U221 ( .A(n211), .B(n206), .Y(n210) );
XOR2X1 U222 ( .A(n212), .B(n213), .Y(N397) );
NOR2X1 U223 ( .A(n214), .B(n198), .Y(n213) );
XOR2X1 U224 ( .A(n215), .B(n216), .Y(N396) );
NOR2X1 U225 ( .A(n217), .B(n198), .Y(n216) );
INVX1 U226 ( .A(G13), .Y(n215) );
XOR2X1 U227 ( .A(n218), .B(n219), .Y(N395) );
NOR2X1 U228 ( .A(n220), .B(n221), .Y(n219) );
XOR2X1 U229 ( .A(n222), .B(n223), .Y(G1355) );
NOR2X1 U230 ( .A(n224), .B(n202), .Y(n223) );
XOR2X1 U231 ( .A(n225), .B(n226), .Y(G1354) );
NOR2X1 U232 ( .A(n205), .B(n202), .Y(n226) );
INVX1 U233 ( .A(n227), .Y(G1352) );
XOR2X1 U234 ( .A(G29), .B(n228), .Y(n227) );
NOR2X1 U235 ( .A(n211), .B(n202), .Y(n228) );
NAND4X1 U236 ( .A(n217), .B(n197), .C(n229), .D(n230), .Y(n202) );
NOR2X1 U237 ( .A(n231), .B(n220), .Y(n229) );
XOR2X1 U238 ( .A(n232), .B(n233), .Y(G1351) );
NOR2X1 U239 ( .A(n224), .B(n234), .Y(n233) );
XOR2X1 U240 ( .A(n235), .B(n236), .Y(G1350) );
NOR2X1 U241 ( .A(n205), .B(n234), .Y(n236) );
INVX1 U242 ( .A(n237), .Y(G1349z) );
XOR2X1 U243 ( .A(G26), .B(n238), .Y(n237) );
NOR2X1 U244 ( .A(n201), .B(n234), .Y(n238) );
XOR2X1 U245 ( .A(n239), .B(n240), .Y(G1348) );
NOR2X1 U246 ( .A(n211), .B(n234), .Y(n240) );
NAND4X1 U247 ( .A(n220), .B(n241), .C(n217), .D(n242), .Y(n234) );
INVX1 U248 ( .A(G25), .Y(n239) );
XOR2X1 U249 ( .A(n243), .B(n244), .Y(G1347) );
XOR2X1 U250 ( .A(keyIn[7]), .B(n245), .Y(n244) );
NOR2X1 U251 ( .A(n224), .B(n206), .Y(n245z) );
NAND4X1 U252 ( .A(n197), .B(n246), .C(n214), .D(n242), .Y(n206) );
INVX1 U253 ( .A(n247), .Y(G1343) );
XOR2X1 U254 ( .A(n248), .B(n249), .Y(n247) );
NOR2X1 U255 ( .A(n224), .B(n250), .Y(n249) );
XOR2X1 U256 ( .A(G20), .B(keyIn[1]), .Y(n248) );
INVX1 U257 ( .A(n251), .Y(G1342) );
XOR2X1 U258 ( .A(G19), .B(n252), .Y(n251) );
NOR2X1 U259 ( .A(n205), .B(n250), .Y(n252) );
XOR2X1 U260 ( .A(n253), .B(n254), .Y(G1341) );
NOR2X1 U261 ( .A(n201), .B(n250), .Y(n254) );
XOR2X1 U262 ( .A(n255), .B(n256), .Y(G1340) );
NOR2X1 U263 ( .A(n211), .B(n250), .Y(n256) );
NAND4X1 U264 ( .A(n214), .B(n220), .C(n257), .D(n258), .Y(n250) );
NOR2X1 U265 ( .A(n231), .B(n217), .Y(n257) );
INVX1 U266 ( .A(n242), .Y(n231) );
OAI33X1 U267 ( .A0(n259), .A1(n260), .A2(n261), .B0(n262), .B1(n263), .B2(n264), .Y(n242) );
INVX1 U268 ( .A(n201), .Y(n262) );
XOR2X1 U269 ( .A(n265), .B(n266), .Y(G1339) );
NOR2X1 U270 ( .A(n220), .B(n198), .Y(n266) );
NAND4X1 U271 ( .A(n211), .B(n261), .C(n267), .D(n205), .Y(n198) );
NOR2X1 U272 ( .A(n268), .B(n201), .Y(n267) );
XOR2X1 U273 ( .A(n269), .B(keyIn[5]), .Y(n265) );
INVX1 U274 ( .A(G16), .Y(n269) );
XOR2X1 U275 ( .A(n270), .B(n271), .Y(G1334) );
NOR2X1 U276 ( .A(n197), .B(n221), .Y(n271) );
INVX1 U277 ( .A(n272), .Y(G1333) );
XOR2X1 U278 ( .A(G10), .B(n273), .Y(n272) );
NOR2X1 U279 ( .A(n214), .B(n221), .Y(n273) );
INVX1 U280 ( .A(n274), .Y(G1332) );
XOR2X1 U281 ( .A(G9), .B(n275), .Y(n274) );
NOR2X1 U282 ( .A(n217), .B(n221), .Y(n275) );
NAND4X1 U283 ( .A(n211), .B(n260), .C(n224), .D(n276), .Y(n221) );
NOR2X1 U284 ( .A(n201), .B(n205), .Y(n260) );
XOR2X1 U285 ( .A(n277), .B(n278), .Y(G1331) );
NOR2X1 U286 ( .A(n220), .B(n279), .Y(n278) );
INVX1 U287 ( .A(G8), .Y(n277) );
XOR2X1 U288 ( .A(n280), .B(n281), .Y(G1330) );
NOR2X1 U289 ( .A(n197), .B(n279), .Y(n281) );
INVX1 U290 ( .A(G7), .Y(n280) );
INVX1 U291 ( .A(n282), .Y(G1329) );
XOR2X1 U292 ( .A(G6), .B(n283), .Y(n282) );
NOR2X1 U293 ( .A(n214), .B(n279), .Y(n283) );
INVX1 U294 ( .A(n284), .Y(G1328) );
XOR2X1 U295 ( .A(n285), .B(n286), .Y(n284) );
NOR2X1 U296 ( .A(n217), .B(n279), .Y(n286) );
NAND4X1 U297 ( .A(n201), .B(n263), .C(n205), .D(n276), .Y(n279) );
NOR2X1 U298 ( .A(n224), .B(n211), .Y(n263) );
XOR2X1 U299 ( .A(n287), .B(n288), .Y(G1327) );
NOR2X1 U300 ( .A(n220), .B(n289), .Y(n288) );
XOR2X1 U301 ( .A(n290), .B(n291), .Y(G1326) );
NOR2X1 U302 ( .A(n197), .B(n289), .Y(n291) );
XOR2X1 U303 ( .A(n292), .B(n293), .Y(G1325) );
NOR2X1 U304 ( .A(n214), .B(n289), .Y(n293) );
XOR2X1 U305 ( .A(n294), .B(n295), .Y(G1324) );
NOR2X1 U306 ( .A(n217), .B(n289), .Y(n295) );
NAND4X1 U307 ( .A(n201), .B(n264), .C(n296), .D(n224), .Y(n289) );
INVX1 U308 ( .A(n261), .Y(n224) );
XOR2X1 U309 ( .A(n297), .B(n298), .Y(n261) );
XOR2X1 U310 ( .A(n299), .B(n300), .Y(n298) );
XOR2X1 U311 ( .A(n243), .B(n301), .Y(n300) );
XOR2X1 U312 ( .A(G24), .B(keyIn[3]), .Y(n243) );
XOR2X1 U313 ( .A(n302), .B(n303), .Y(n299) );
NAND2X1 U314 ( .A(G40), .B(G41), .Y(n302) );
XOR2X1 U315 ( .A(n304), .B(n305), .Y(n297) );
XOR2X1 U316 ( .A(keyIn[4]), .B(G32), .Y(n305) );
XOR2X1 U317 ( .A(G20), .B(n232), .Y(n304) );
NOR2X1 U318 ( .A(n268), .B(n211), .Y(n296) );
INVX1 U319 ( .A(n259), .Y(n211) );
XOR2X1 U320 ( .A(n306), .B(n307), .Y(n259) );
XOR2X1 U321 ( .A(n308), .B(n309), .Y(n307) );
XOR2X1 U322 ( .A(n310), .B(n301), .Y(n309) );
XOR2X1 U323 ( .A(n311), .B(n312), .Y(n301) );
XOR2X1 U324 ( .A(G6), .B(n285), .Y(n312) );
XOR2X1 U325 ( .A(G5), .B(keyIn[6]), .Y(n285) );
XOR2X1 U326 ( .A(G7), .B(G8), .Y(n311) );
XOR2X1 U327 ( .A(n255), .B(n313), .Y(n308) );
NAND2X1 U328 ( .A(G37), .B(G41), .Y(n313) );
XOR2X1 U329 ( .A(n314), .B(n315), .Y(n306) );
XOR2X1 U330 ( .A(keyIn[0]), .B(G29), .Y(n315) );
XOR2X1 U331 ( .A(n209), .B(G25), .Y(n314) );
INVX1 U332 ( .A(G21), .Y(n209) );
INVX1 U333 ( .A(n276), .Y(n268) );
OAI33X1 U334 ( .A0(n316), .A1(n241), .A2(n317), .B0(n258), .B1(n246), .B2(n230), .Y(n276) );
INVX1 U335 ( .A(n214), .Y(n230) );
NOR2X1 U336 ( .A(n217), .B(n220), .Y(n246) );
INVX1 U337 ( .A(n316), .Y(n220) );
INVX1 U338 ( .A(n197), .Y(n258) );
NOR2X1 U339 ( .A(n214), .B(n197), .Y(n241) );
XOR2X1 U340 ( .A(n318), .B(n319), .Y(n197) );
XOR2X1 U341 ( .A(n320), .B(n321), .Y(n319) );
XOR2X1 U342 ( .A(n322), .B(n323), .Y(n321) );
NAND2X1 U343 ( .A(G35), .B(G41), .Y(n322) );
XOR2X1 U344 ( .A(n324), .B(n325), .Y(n318) );
XOR2X1 U345 ( .A(G7), .B(G3), .Y(n325) );
XOR2X1 U346 ( .A(n270), .B(G15), .Y(n324) );
INVX1 U347 ( .A(G11), .Y(n270) );
XOR2X1 U348 ( .A(n326), .B(n327), .Y(n214) );
XOR2X1 U349 ( .A(n328), .B(n329), .Y(n327) );
XOR2X1 U350 ( .A(n330), .B(n323), .Y(n329) );
XOR2X1 U351 ( .A(n331), .B(n332), .Y(n323) );
XOR2X1 U352 ( .A(n232), .B(n235), .Y(n332) );
INVX1 U353 ( .A(G28), .Y(n232) );
XOR2X1 U354 ( .A(G25), .B(G26), .Y(n331) );
NAND2X1 U355 ( .A(G34), .B(G41), .Y(n330z) );
XOR2X1 U356 ( .A(n333), .B(n334), .Y(n326) );
XOR2X1 U357 ( .A(G6), .B(G2), .Y(n334) );
XOR2X1 U358 ( .A(G10), .B(n212), .Y(n333) );
XOR2X1 U359 ( .A(n335), .B(n336), .Y(n316) );
XOR2X1 U360 ( .A(n328), .B(n337), .Y(n336) );
XOR2X1 U361 ( .A(n338), .B(n339), .Y(n337) );
NAND2X1 U362 ( .A(G41), .B(G36), .Y(n338) );
XOR2X1 U363 ( .A(n340), .B(n341), .Y(n328) );
XOR2X1 U364 ( .A(n222), .B(n225), .Y(n341) );
INVX1 U365 ( .A(G32), .Y(n222) );
XOR2X1 U366 ( .A(G29), .B(n199), .Y(n340) );
INVX1 U367 ( .A(G30), .Y(n199) );
XOR2X1 U368 ( .A(n342), .B(n343), .Y(n335) );
XOR2X1 U369 ( .A(G8), .B(G4), .Y(n343) );
XOR2X1 U370 ( .A(n218), .B(G16), .Y(n342) );
INVX1 U371 ( .A(G12), .Y(n218) );
INVX1 U372 ( .A(n205), .Y(n264) );
XOR2X1 U373 ( .A(n344), .B(n345), .Y(n205) );
XOR2X1 U374 ( .A(n310), .B(n346), .Y(n345) );
XOR2X1 U375 ( .A(n347), .B(n348), .Y(n346) );
NAND2X1 U376 ( .A(G39), .B(G41), .Y(n347) );
XOR2X1 U377 ( .A(n349), .B(n350), .Y(n310) );
XOR2X1 U378 ( .A(n287), .B(n290), .Y(n350) );
INVX1 U379 ( .A(G3), .Y(n290) );
INVX1 U380 ( .A(G4), .Y(n287) );
XOR2X1 U381 ( .A(G1), .B(n292), .Y(n349) );
INVX1 U382 ( .A(G2), .Y(n292z) );
XOR2X1 U383 ( .A(n351), .B(n352), .Y(n344) );
XOR2X1 U384 ( .A(n225), .B(n235), .Y(n352z) );
INVX1 U385 ( .A(G27), .Y(n235) );
INVX1 U386 ( .A(G31), .Y(n225) );
XOR2X1 U387 ( .A(G19), .B(n203), .Y(n351) );
INVX1 U388 ( .A(G23), .Y(n203) );
XOR2X1 U389 ( .A(n353), .B(n354), .Y(n201) );
XOR2X1 U390 ( .A(n303), .B(n355), .Y(n354) );
XOR2X1 U391 ( .A(n356), .B(n348), .Y(n355) );
XOR2X1 U392 ( .A(n357), .B(n358), .Y(n348) );
XOR2X1 U393 ( .A(G9), .B(G12), .Y(n358) );
XOR2X1 U394 ( .A(G10), .B(G11), .Y(n357) );
NAND2X1 U395 ( .A(G38), .B(G41), .Y(n356) );
XOR2X1 U396 ( .A(n359), .B(n360), .Y(n303) );
XOR2X1 U397 ( .A(G16), .B(G15), .Y(n360) );
XOR2X1 U398 ( .A(G13), .B(n212), .Y(n359) );
INVX1 U399 ( .A(G14), .Y(n212) );
XOR2X1 U400 ( .A(n361), .B(n362), .Y(n353) );
XOR2X1 U401 ( .A(G30), .B(G26), .Y(n362) );
XOR2X1 U402 ( .A(n253), .B(G22), .Y(n361) );
INVX1 U403 ( .A(G18), .Y(n253) );
INVX1 U404 ( .A(n317), .Y(n217) );
XOR2X1 U405 ( .A(n363), .B(n364), .Y(n317) );
XOR2X1 U406 ( .A(n339), .B(n365), .Y(n364) );
XOR2X1 U407 ( .A(n366), .B(n320), .Y(n365z) );
XOR2X1 U408 ( .A(n367), .B(n368), .Y(n320z) );
XOR2X1 U409 ( .A(G20), .B(G19), .Y(n368) );
XOR2X1 U410 ( .A(n255), .B(G18), .Y(n367) );
INVX1 U411 ( .A(G17), .Y(n255) );
NAND2X1 U412 ( .A(G33), .B(G41), .Y(n366) );
XOR2X1 U413 ( .A(n369), .B(n370), .Y(n339) );
XOR2X1 U414 ( .A(G24), .B(G23), .Y(n370z) );
XOR2X1 U415 ( .A(G21), .B(n207), .Y(n369) );
INVX1 U416 ( .A(G22), .Y(n207) );
XOR2X1 U417 ( .A(n371), .B(n372), .Y(n363) );
XOR2X1 U418 ( .A(G9), .B(G5), .Y(n372) );
XOR2X1 U419 ( .A(n294), .B(G13), .Y(n371) );
INVX1 U420 ( .A(G1), .Y(n294) );
  XOR2X1 enc2XOR2X10 ( .A(keyInPseudo[2]), .B(n365z), .Y(n365z_inv_wire) );
  INVX1 inv0inv( .A(n365z_inv_wire), .Y(n365) );
  XOR2X1 enc2XOR2X11 ( .A(keyInPseudo[6]), .B(n352z), .Y(n352z_inv_wire) );
  INVX1 inv1inv( .A(n352z_inv_wire), .Y(n352) );
  XOR2X1 enc2XOR2X12 ( .A(keyInPseudo[5]), .B(G1349z), .Y(G1349) );
  XOR2X1 enc2XOR2X13 ( .A(keyInPseudo[3]), .B(n245z), .Y(n245) );
  XOR2X1 enc2XOR2X14 ( .A(keyInPseudo[4]), .B(n370z), .Y(n370) );
  XOR2X1 enc2XOR2X15 ( .A(keyInPseudo[0]), .B(n330z), .Y(n330z_inv_wire) );
  INVX1 inv2inv( .A(n330z_inv_wire), .Y(n330) );
  XOR2X1 enc2XOR2X16 ( .A(keyInPseudo[1]), .B(n320z), .Y(n320) );
  XOR2X1 enc2XOR2X17 ( .A(keyInPseudo[7]), .B(n292z), .Y(n292) );
endmodule