// keyIn= 10001111
module c1355 (keyIn,  G1,  G10,  G11,  G12,  G13,  G14,  G15,  G16,  G17,  G18,  G19,  G2,  G20,  G21,  G22,  G23,  G24,  G25,  G26,  G27,  G28,  G29,  G3,  G30,  G31,  G32,  G33,  G34,  G35,  G36,  G37,  G38,  G39,  G4,  G40,  G41,  G5,  G6,  G7,  G8,  G9,  G1324,  G1325,  G1326,  G1327,  G1328,  G1329,  G1330,  G1331,  G1332,  G1333,  G1334,  G1335,  G1336,  G1337,  G1338,  G1339,  G1340,  G1341,  G1342,  G1343,  G1344,  G1345,  G1346,  G1347,  G1348,  G1349,  G1350,  G1351,  G1352,  G1353,  G1354,  G1355 ); 
input [7:0] keyIn; 
input G1, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9; 
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355; 
wire   N388, N395, N396, N397, N404, N405, N406, N407, N409, N413, n17678, n17679, n17680, n17681, n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689, n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697, n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705, n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713, n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721, n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729, n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737, n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745, n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753, n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761, n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769, n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777, n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785, n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793, n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801, n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809, n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817, n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825, n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833, n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841, n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849; 
assign G1328 = N388;
assign G1335 = N395;
assign G1336 = N396;
assign G1337 = N397;
assign G1344 = N404;
assign G1345 = N405;
assign G1346 = N406;
assign G1347 = N407;
assign G1349 = N409;
assign G1353 = N413;
XOR2X1 U10281 ( .A(n17678), .B(n17679), .Y(N413) );
NOR2X1 U10282 ( .A(n17680), .B(n17681), .Y(n17679) );
XOR2X1 U10283 ( .A(n17682), .B(n17683), .Y(N409) );
NOR2X1 U10284 ( .A(n17680), .B(n17684), .Y(n17683) );
XOR2X1 U10285 ( .A(n17685), .B(n17686), .Y(N407) );
NOR2X1 U10286 ( .A(n17687), .B(n17688), .Y(n17686) );
XOR2X1 U10287 ( .A(n17689), .B(n17690), .Y(N406) );
NOR2X1 U10288 ( .A(n17691), .B(n17688), .Y(n17690) );
XOR2X1 U10289 ( .A(n17692), .B(n17693), .Y(N405) );
NOR2X1 U10290 ( .A(n17680), .B(n17688), .Y(n17693) );
XOR2X1 U10291 ( .A(n17694), .B(n17695), .Y(N404) );
NOR2X1 U10292 ( .A(n17696), .B(n17688), .Y(n17695) );
NAND4X1 U10293 ( .A(n17697), .B(n17698), .C(n17699), .D(n17700), .Y(n17688) );
NOR2X1 U10294 ( .A(n17701), .B(n17702), .Y(n17699) );
XOR2X1 U10295 ( .A(n17703), .B(n17704), .Y(N397) );
NOR2X1 U10296 ( .A(n17697), .B(n17705), .Y(n17704) );
XOR2X1 U10297 ( .A(n17706), .B(n17707), .Y(N396) );
NOR2X1 U10298 ( .A(n17708), .B(n17705), .Y(n17707) );
XOR2X1 U10299 ( .A(n17709), .B(n17710), .Y(N395) );
NOR2X1 U10300 ( .A(n17702), .B(n17711), .Y(n17710) );
XOR2X1 U10301 ( .A(n17712), .B(n17713), .Y(N388) );
NOR2X1 U10302 ( .A(n17708), .B(n17714), .Y(n17713) );
INVX1 U10303 ( .A(n17715), .Y(G1355) );
XOR2X1 U10304 ( .A(G32), .B(n17716), .Y(n17715) );
NOR2X1 U10305 ( .A(n17687), .B(n17681), .Y(n17716) );
INVX1 U10306 ( .A(n17717), .Y(G1354) );
XOR2X1 U10307 ( .A(G31), .B(n17718), .Y(n17717z) );
NOR2X1 U10308 ( .A(n17691), .B(n17681), .Y(n17718) );
XOR2X1 U10309 ( .A(n17719), .B(n17720), .Y(G1352) );
NOR2X1 U10310 ( .A(n17696), .B(n17681), .Y(n17720) );
NAND4X1 U10311 ( .A(n17698), .B(n17721), .C(n17708), .D(n17722), .Y(n17681) );
INVX1 U10312 ( .A(G29), .Y(n17719) );
INVX1 U10313 ( .A(n17723), .Y(G1351) );
XOR2X1 U10314 ( .A(G28), .B(n17724), .Y(n17723) );
NOR2X1 U10315 ( .A(n17687), .B(n17684), .Y(n17724) );
INVX1 U10316 ( .A(n17725), .Y(G1350) );
XOR2X1 U10317 ( .A(G27), .B(n17726), .Y(n17725) );
NOR2X1 U10318 ( .A(n17691), .B(n17684), .Y(n17726) );
XOR2X1 U10319 ( .A(n17727), .B(n17728), .Y(G1348) );
NOR2X1 U10320 ( .A(n17696), .B(n17684), .Y(n17728) );
NAND4X1 U10321 ( .A(n17702), .B(n17708), .C(n17729), .D(n17730), .Y(n17684z) );
NOR2X1 U10322 ( .A(n17701), .B(n17697), .Y(n17729) );
INVX1 U10323 ( .A(n17722), .Y(n17701) );
INVX1 U10324 ( .A(G25), .Y(n17727) );
XOR2X1 U10325 ( .A(n17731), .B(n17732), .Y(G1343) );
NOR2X1 U10326 ( .A(n17687), .B(n17733), .Y(n17732) );
INVX1 U10327 ( .A(G20), .Y(n17731) );
XOR2X1 U10328 ( .A(n17734), .B(n17735), .Y(G1342) );
NOR2X1 U10329 ( .A(n17691), .B(n17733), .Y(n17735) );
INVX1 U10330 ( .A(G19), .Y(n17734) );
XOR2X1 U10331 ( .A(n17736), .B(n17737), .Y(G1341) );
NOR2X1 U10332 ( .A(n17680), .B(n17733), .Y(n17737) );
INVX1 U10333 ( .A(G18), .Y(n17736) );
XOR2X1 U10334 ( .A(n17738), .B(n17739), .Y(G1340) );
NOR2X1 U10335 ( .A(n17696), .B(n17733), .Y(n17739) );
NAND4X1 U10336 ( .A(n17697), .B(n17740), .C(n17702), .D(n17722), .Y(n17733) );
OAI33X1 U10337 ( .A0(n17741), .A1(n17742), .A2(n17743), .B0(n17744), .B1(n17745), .B2(n17746), .Y(n17722) );
INVX1 U10338 ( .A(n17696), .Y(n17743) );
INVX1 U10339 ( .A(n17691), .Y(n17741) );
INVX1 U10340 ( .A(G17), .Y(n17738) );
INVX1 U10341 ( .A(n17747), .Y(G1339) );
XOR2X1 U10342 ( .A(G16), .B(n17748), .Y(n17747) );
NOR2X1 U10343 ( .A(n17702), .B(n17705), .Y(n17748) );
INVX1 U10344 ( .A(n17749), .Y(G1338) );
XOR2X1 U10345 ( .A(G15), .B(n17750), .Y(n17749) );
NOR2X1 U10346 ( .A(n17698), .B(n17705), .Y(n17750) );
NAND4X1 U10347 ( .A(n17691), .B(n17742), .C(n17696), .D(n17751), .Y(n17705) );
NOR2X1 U10348 ( .A(n17687), .B(n17680), .Y(n17742) );
XOR2X1 U10349 ( .A(n17752), .B(n17753), .Y(G1334) );
NOR2X1 U10350 ( .A(n17698), .B(n17711), .Y(n17753) );
XOR2X1 U10351 ( .A(n17754), .B(n17755), .Y(G1333) );
NOR2X1 U10352 ( .A(n17697), .B(n17711), .Y(n17755) );
INVX1 U10353 ( .A(n17756), .Y(G1332) );
XOR2X1 U10354 ( .A(G9), .B(n17757), .Y(n17756) );
NOR2X1 U10355 ( .A(n17708), .B(n17711), .Y(n17757) );
NAND4X1 U10356 ( .A(n17687), .B(n17696), .C(n17758), .D(n17744), .Y(n17711) );
INVX1 U10357 ( .A(n17680), .Y(n17744) );
NOR2X1 U10358 ( .A(n17759), .B(n17691), .Y(n17758) );
INVX1 U10359 ( .A(n17760), .Y(G1331) );
XOR2X1 U10360 ( .A(G8), .B(n17761), .Y(n17760) );
NOR2X1 U10361 ( .A(n17702), .B(n17714), .Y(n17761) );
INVX1 U10362 ( .A(n17762), .Y(G1330) );
XOR2X1 U10363 ( .A(G7), .B(n17763), .Y(n17762) );
NOR2X1 U10364 ( .A(n17698), .B(n17714), .Y(n17763) );
INVX1 U10365 ( .A(n17764), .Y(G1329) );
XOR2X1 U10366 ( .A(G6), .B(n17765), .Y(n17764) );
NOR2X1 U10367 ( .A(n17697), .B(n17714), .Y(n17765) );
NAND4X1 U10368 ( .A(n17691), .B(n17680), .C(n17766), .D(n17746), .Y(n17714z) );
INVX1 U10369 ( .A(n17687), .Y(n17746) );
NOR2X1 U10370 ( .A(n17759), .B(n17696), .Y(n17766) );
INVX1 U10371 ( .A(n17751), .Y(n17759) );
INVX1 U10372 ( .A(n17767), .Y(G1327) );
XOR2X1 U10373 ( .A(G4), .B(n17768), .Y(n17767) );
NOR2X1 U10374 ( .A(n17702), .B(n17769), .Y(n17768) );
INVX1 U10375 ( .A(n17770), .Y(G1326) );
XOR2X1 U10376 ( .A(G3), .B(n17771), .Y(n17770) );
NOR2X1 U10377 ( .A(n17698), .B(n17769), .Y(n17771) );
XOR2X1 U10378 ( .A(n17772), .B(n17773), .Y(G1325) );
NOR2X1 U10379 ( .A(n17697), .B(n17769), .Y(n17773) );
XOR2X1 U10380 ( .A(n17774), .B(n17775), .Y(G1324) );
NOR2X1 U10381 ( .A(n17708), .B(n17769), .Y(n17775z) );
NAND4X1 U10382 ( .A(n17680), .B(n17745), .C(n17687), .D(n17751), .Y(n17769) );
OAI33X1 U10383 ( .A0(n17730), .A1(n17721), .A2(n17700), .B0(n17776), .B1(n17740), .B2(n17777), .Y(n17751) );
NOR2X1 U10384 ( .A(n17708), .B(n17698), .Y(n17740) );
INVX1 U10385 ( .A(n17708), .Y(n17700) );
NOR2X1 U10386 ( .A(n17702), .B(n17697), .Y(n17721) );
INVX1 U10387 ( .A(n17776), .Y(n17697) );
XOR2X1 U10388 ( .A(n17778), .B(n17779), .Y(n17776) );
XOR2X1 U10389 ( .A(n17780), .B(n17781), .Y(n17779) );
XOR2X1 U10390 ( .A(n17782), .B(n17783), .Y(n17781) );
NAND2X1 U10391 ( .A(G34), .B(G41), .Y(n17782z) );
XOR2X1 U10392 ( .A(n17784), .B(n17785), .Y(n17778) );
XOR2X1 U10393 ( .A(G6), .B(G2), .Y(n17785) );
XOR2X1 U10394 ( .A(G10), .B(n17703), .Y(n17784) );
INVX1 U10395 ( .A(n17777), .Y(n17702) );
XOR2X1 U10396 ( .A(n17786), .B(n17787), .Y(n17777z) );
XOR2X1 U10397 ( .A(n17780), .B(n17788), .Y(n17787) );
XOR2X1 U10398 ( .A(n17789), .B(n17790), .Y(n17788) );
NAND2X1 U10399 ( .A(G36), .B(G41), .Y(n17789) );
XOR2X1 U10400 ( .A(n17791), .B(n17792), .Y(n17780) );
XOR2X1 U10401 ( .A(G32), .B(G31), .Y(n17792) );
XOR2X1 U10402 ( .A(G29), .B(n17678), .Y(n17791) );
INVX1 U10403 ( .A(G30), .Y(n17678) );
XOR2X1 U10404 ( .A(n17793), .B(n17794), .Y(n17786) );
XOR2X1 U10405 ( .A(G8), .B(G4), .Y(n17794) );
XOR2X1 U10406 ( .A(n17709), .B(G16), .Y(n17793) );
INVX1 U10407 ( .A(G12), .Y(n17709) );
INVX1 U10408 ( .A(n17698), .Y(n17730) );
XOR2X1 U10409 ( .A(n17795), .B(n17796), .Y(n17698) );
XOR2X1 U10410 ( .A(n17783), .B(n17797), .Y(n17796) );
XOR2X1 U10411 ( .A(n17798), .B(n17799), .Y(n17797) );
NAND2X1 U10412 ( .A(G35), .B(G41), .Y(n17798) );
XOR2X1 U10413 ( .A(n17800), .B(n17801), .Y(n17783) );
XOR2X1 U10414 ( .A(G28), .B(G27), .Y(n17801) );
XOR2X1 U10415 ( .A(G25), .B(n17682), .Y(n17800) );
INVX1 U10416 ( .A(G26), .Y(n17682) );
XOR2X1 U10417 ( .A(n17802), .B(n17803), .Y(n17795) );
XOR2X1 U10418 ( .A(G7), .B(G3), .Y(n17803) );
XOR2X1 U10419 ( .A(n17752), .B(G15), .Y(n17802) );
INVX1 U10420 ( .A(G11), .Y(n17752) );
XOR2X1 U10421 ( .A(n17804), .B(n17805), .Y(n17687) );
XOR2X1 U10422 ( .A(n17806), .B(n17807), .Y(n17805) );
XOR2X1 U10423 ( .A(n17808), .B(n17809), .Y(n17807) );
NAND2X1 U10424 ( .A(G40), .B(G41), .Y(n17808) );
XOR2X1 U10425 ( .A(n17810), .B(n17811), .Y(n17804) );
XOR2X1 U10426 ( .A(G32), .B(G28), .Y(n17811) );
XOR2X1 U10427 ( .A(G20), .B(n17685), .Y(n17810) );
INVX1 U10428 ( .A(G24), .Y(n17685) );
NOR2X1 U10429 ( .A(n17696), .B(n17691), .Y(n17745) );
XOR2X1 U10430 ( .A(n17812), .B(n17813), .Y(n17691) );
XOR2X1 U10431 ( .A(n17814), .B(n17815), .Y(n17813) );
XOR2X1 U10432 ( .A(n17816), .B(n17817), .Y(n17815) );
NAND2X1 U10433 ( .A(G41), .B(G39), .Y(n17816) );
XOR2X1 U10434 ( .A(n17818), .B(n17819), .Y(n17812) );
XOR2X1 U10435 ( .A(G31), .B(G27), .Y(n17819) );
XOR2X1 U10436 ( .A(G19), .B(n17689), .Y(n17818) );
INVX1 U10437 ( .A(G23), .Y(n17689) );
XOR2X1 U10438 ( .A(n17820), .B(n17821), .Y(n17696) );
XOR2X1 U10439 ( .A(n17806), .B(n17822), .Y(n17821) );
XOR2X1 U10440 ( .A(n17823), .B(n17814), .Y(n17822) );
XOR2X1 U10441 ( .A(n17824), .B(n17825), .Y(n17814) );
XOR2X1 U10442 ( .A(G4), .B(G3), .Y(n17825) );
XOR2X1 U10443 ( .A(n17774), .B(n17772), .Y(n17824) );
INVX1 U10444 ( .A(G2), .Y(n17772) );
NAND2X1 U10445 ( .A(G37), .B(G41), .Y(n17823) );
XOR2X1 U10446 ( .A(n17826), .B(n17827), .Y(n17806) );
XOR2X1 U10447 ( .A(G8), .B(G7), .Y(n17827) );
XOR2X1 U10448 ( .A(n17712), .B(G6), .Y(n17826) );
INVX1 U10449 ( .A(G5), .Y(n17712) );
XOR2X1 U10450 ( .A(n17828), .B(n17829), .Y(n17820) );
XOR2X1 U10451 ( .A(G29), .B(G25), .Y(n17829z) );
XOR2X1 U10452 ( .A(G17), .B(n17694), .Y(n17828) );
XOR2X1 U10453 ( .A(n17830), .B(n17831), .Y(n17680) );
XOR2X1 U10454 ( .A(n17817), .B(n17832), .Y(n17831) );
XOR2X1 U10455 ( .A(n17833), .B(n17809), .Y(n17832z) );
XOR2X1 U10456 ( .A(n17834), .B(n17835), .Y(n17809) );
XOR2X1 U10457 ( .A(G16), .B(G15), .Y(n17835) );
XOR2X1 U10458 ( .A(n17706), .B(n17703), .Y(n17834) );
INVX1 U10459 ( .A(G14), .Y(n17703) );
NAND2X1 U10460 ( .A(G38), .B(G41), .Y(n17833) );
XOR2X1 U10461 ( .A(n17836), .B(n17837), .Y(n17817) );
XOR2X1 U10462 ( .A(G9), .B(G12), .Y(n17837) );
XOR2X1 U10463 ( .A(n17754), .B(G11), .Y(n17836) );
INVX1 U10464 ( .A(G10), .Y(n17754) );
XOR2X1 U10465 ( .A(n17838), .B(n17839), .Y(n17830) );
XOR2X1 U10466 ( .A(G30), .B(G26), .Y(n17839) );
XOR2X1 U10467 ( .A(G18), .B(n17692), .Y(n17838) );
INVX1 U10468 ( .A(G22), .Y(n17692) );
XOR2X1 U10469 ( .A(n17840), .B(n17841), .Y(n17708) );
XOR2X1 U10470 ( .A(n17790), .B(n17842), .Y(n17841) );
XOR2X1 U10471 ( .A(n17843), .B(n17799), .Y(n17842) );
XOR2X1 U10472 ( .A(n17844), .B(n17845), .Y(n17799) );
XOR2X1 U10473 ( .A(G20), .B(G19), .Y(n17845) );
XOR2X1 U10474 ( .A(G17), .B(G18), .Y(n17844) );
NAND2X1 U10475 ( .A(G33), .B(G41), .Y(n17843) );
XOR2X1 U10476 ( .A(n17846), .B(n17847), .Y(n17790) );
XOR2X1 U10477 ( .A(G24), .B(G23), .Y(n17847) );
XOR2X1 U10478 ( .A(n17694), .B(G22), .Y(n17846) );
INVX1 U10479 ( .A(G21), .Y(n17694) );
XOR2X1 U10480 ( .A(n17848), .B(n17849), .Y(n17840) );
XOR2X1 U10481 ( .A(G9), .B(G5), .Y(n17849) );
XOR2X1 U10482 ( .A(G1), .B(n17706), .Y(n17848) );
INVX1 U10483 ( .A(G13), .Y(n17706) );
INVX1 U10484 ( .A(G1), .Y(n17774) );
  XOR2X1 encXOR2X10 ( .A(n17684z), .B(keyIn[7]), .Y(n17684z_inv_wire) );
  INVX1 encgate0inv( .A(n17684z_inv_wire), .Y(n17684) );
  XOR2X1 encXOR2X11 ( .A(keyIn[2]), .B(n17777z), .Y(n17777) );
  XOR2X1 encXOR2X12 ( .A(n17782z), .B(keyIn[4]), .Y(n17782z_inv_wire) );
  INVX1 encgate2inv( .A(n17782z_inv_wire), .Y(n17782) );
  XOR2X1 encXOR2X13 ( .A(n17717z), .B(keyIn[6]), .Y(n17717z_inv_wire) );
  INVX1 encgate3inv( .A(n17717z_inv_wire), .Y(n17717) );
  XOR2X1 encXOR2X14 ( .A(keyIn[1]), .B(n17714z), .Y(n17714) );
  XOR2X1 encXOR2X15 ( .A(n17829z), .B(keyIn[5]), .Y(n17829z_inv_wire) );
  INVX1 encgate5inv( .A(n17829z_inv_wire), .Y(n17829) );
  XOR2X1 encXOR2X16 ( .A(keyIn[3]), .B(n17832z), .Y(n17832) );
  XOR2X1 encXOR2X17 ( .A(n17775z), .B(keyIn[0]), .Y(n17775z_inv_wire) );
  INVX1 encgate7inv( .A(n17775z_inv_wire), .Y(n17775) );
endmodule