// key= 10000010
module c2670 (keyInPseudo,  keyIn,  G1,  G10,  G100,  G101,  G102,  G103,  G104,  G105,  G106,  G107,  G108,  G109,  G11,  G110,  G111,  G112,  G113,  G114,  G115,  G116,  G117,  G118,  G119,  G12,  G120,  G121,  G122,  G123,  G124,  G125,  G126,  G127,  G128,  G129,  G13,  G130,  G131,  G132,  G133,  G134,  G135,  G136,  G137,  G138,  G139,  G14,  G140,  G141,  G142,  G143,  G144,  G145,  G146,  G147,  G148,  G149,  G15,  G150,  G151,  G152,  G153,  G154,  G155,  G156,  G157,  G16,  G17,  G18,  G19,  G2,  G20,  G21,  G22,  G23,  G24,  G25,  G26,  G27,  G28,  G29,  G3,  G30,  G31,  G32,  G33,  G34,  G35,  G36,  G37,  G38,  G39,  G4,  G40,  G41,  G42,  G43,  G44,  G45,  G46,  G47,  G48,  G49,  G5,  G50,  G51,  G52,  G53,  G54,  G55,  G56,  G57,  G58,  G59,  G6,  G60,  G61,  G62,  G63,  G64,  G65,  G66,  G67,  G68,  G69,  G7,  G70,  G71,  G72,  G73,  G74,  G75,  G76,  G77,  G78,  G79,  G8,  G80,  G81,  G82,  G83,  G84,  G85,  G86,  G87,  G88,  G89,  G9,  G90,  G91,  G92,  G93,  G94,  G95,  G96,  G97,  G98,  G99,  G2531,  G2532,  G2533,  G2534,  G2535,  G2536,  G2537,  G2538,  G2539,  G2540,  G2541,  G2542,  G2543,  G2544,  G2545,  G2546,  G2547,  G2548,  G2549,  G2550,  G2551,  G2552,  G2553,  G2554,  G2555,  G2556,  G2557,  G2558,  G2559,  G2560,  G2561,  G2562,  G2563,  G2564,  G2565,  G2566,  G2567,  G2568,  G2569,  G2570,  G2571,  G2572,  G2573,  G2574,  G2575,  G2576,  G2577,  G2578,  G2579,  G2580,  G2581,  G2582,  G2583,  G2584,  G2585,  G2586,  G2587,  G2588,  G2589,  G2590,  G2591,  G2592,  G2593,  G2594 ); 
input [7:0] keyIn; 
input  [7:0] keyInPseudo; 
input G1, G10, G100, G101, G102, G103, G104, G105, G106, G107, G108, G109, G11, G110, G111, G112, G113, G114, G115, G116, G117, G118, G119, G12, G120, G121, G122, G123, G124, G125, G126, G127, G128, G129, G13, G130, G131, G132, G133, G134, G135, G136, G137, G138, G139, G14, G140, G141, G142, G143, G144, G145, G146, G147, G148, G149, G15, G150, G151, G152, G153, G154, G155, G156, G157, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G42, G43, G44, G45, G46, G47, G48, G49, G5, G50, G51, G52, G53, G54, G55, G56, G57, G58, G59, G6, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G7, G70, G71, G72, G73, G74, G75, G76, G77, G78, G79, G8, G80, G81, G82, G83, G84, G85, G86, G87, G88, G89, G9, G90, G91, G92, G93, G94, G95, G96, G97, G98, G99; 
output G2531, G2532, G2533, G2534, G2535, G2536, G2537, G2538, G2539, G2540, G2541, G2542, G2543, G2544, G2545, G2546, G2547, G2548, G2549, G2550, G2551, G2552, G2553, G2554, G2555, G2556, G2557, G2558, G2559, G2560, G2561, G2562, G2563, G2564, G2565, G2566, G2567, G2568, G2569, G2570, G2571, G2572, G2573, G2574, G2575, G2576, G2577, G2578, G2579, G2580, G2581, G2582, G2583, G2584, G2585, G2586, G2587, G2588, G2589, G2590, G2591, G2592, G2593, G2594; 
wire   N155, G115, G1014, G1017, G1021, G1026, G1030, G1033, G1036, G2594, G2585, G2555, G2531, G2589, G2576, G2574, G2579, G2534, G2536, n25076, n25077, n25078, n25079, n25080, n25081, n25082, n25083, n25084, n25085, n25086, n25087, n25088, n25089, n25090, n25091, n25092, n25093, n25094, n25095, n25096, n25097, n25098, n25099, n25100, n25101, n25102, n25103, n25104, n25105, n25106, n25107, n25108, n25109, n25110, n25111, n25112, n25113, n25114, n25115, n25116, n25117, n25118, n25119, n25120, n25121, n25122, n25123, n25124, n25125, n25126, n25127, n25128, n25129, n25130, n25131, n25132, n25133, n25134, n25135, n25136, n25137, n25138, n25139, n25140, n25141, n25142, n25143, n25144, n25145, n25146, n25147, n25148, n25149, n25150, n25151, n25152, n25153, n25154, n25155, n25156, n25157, n25158, n25159, n25160, n25161, n25162, n25163, n25164, n25165, n25166, n25167, n25168, n25169, n25170, n25171, n25172, n25173, n25174, n25175, n25176, n25177, n25178, n25179, n25180, n25181, n25182, n25183, n25184, n25185, n25186, n25187, n25188, n25189, n25190, n25191, n25192, n25193, n25194, n25195, n25196, n25197, n25198, n25199, n25200, n25201, n25202, n25203, n25204, n25205, n25206, n25207, n25208, n25209, n25210, n25211, n25212, n25213, n25214, n25215, n25216, n25217, n25218, n25219, n25220, n25221, n25222, n25223, n25224, n25225, n25226, n25227, n25228, n25229, n25230, n25231, n25232, n25233, n25234, n25235, n25236, n25237, n25238, n25239, n25240, n25241, n25242, n25243, n25244, n25245, n25246, n25247, n25248, n25249, n25250, n25251, n25252, n25253, n25254, n25255, n25256, n25257, n25258, n25259, n25260, n25261, n25262, n25263, n25264, n25265, n25266, n25267, n25268, n25269, n25270, n25271, n25272, n25273, n25274, n25275, n25276, n25277, n25278, n25279, n25280, n25281, n25282, n25283, n25284, n25285, n25286, n25287, n25288, n25289, n25290, n25291, n25292, n25293, n25294, n25295, n25296, n25297, n25298, n25299, n25300, n25301, n25302, n25303, n25304, n25305, n25306, n25307, n25308, n25309, n25310, n25311, n25312; 
assign G2549 = G115;
assign G2554 = G2555;
assign G2584 = G2585;
assign G2592 = 1'b0;
assign G2593 = G2594;
assign G2582 = N155;
assign G2566 = G1014;
assign G2567 = G1017;
assign G2568 = G1021;
assign G2569z = G1026;
assign G2570 = G1030;
assign G2571 = G1033;
assign G2572 = G1036;
assign G2588 = G2589;
assign G2575 = G2576;
assign G2533z = G2531;
assign G2532 = G2531;
assign G2573 = G2574;
assign G2578 = G2579;
assign G2535 = G2534;
assign G2536 = G2538;
assign G2537 = G2538;
NAND4X1 U301 ( .A(G2590), .B(n273), .C(G2587), .D(n274), .Y(G2594) );
NOR2X1 U302 ( .A(G2583), .B(n275), .Y(n274) );
NAND2X1 U303 ( .A(n276), .B(G2581), .Y(n275) );
INVX1 U304 ( .A(N155), .Y(n276) );
XOR2X1 U305 ( .A(n277), .B(n278), .Y(N155) );
XOR2X1 U306 ( .A(n279), .B(n280), .Y(n278) );
XOR2X1 U307 ( .A(G139), .B(G138), .Y(n280) );
XOR2X1 U308 ( .A(G141), .B(G140), .Y(n279) );
XOR2X1 U309 ( .A(n281), .B(n282), .Y(n277) );
XOR2X1 U310 ( .A(G157), .B(G144), .Y(n282) );
XOR2X1 U311 ( .A(G143), .B(n283), .Y(n281) );
AOI21X1 U312 ( .A0(n284), .A1(n285), .B0(n286), .Y(G2591) );
OAI21X1 U313 ( .A0(n287), .A1(n288), .B0(n289), .Y(n286) );
NAND3X1 U314 ( .A(n290), .B(n291), .C(n292), .Y(n289) );
INVX1 U315 ( .A(n293), .Y(n292) );
AOI21X1 U316 ( .A0(n294), .A1(n285), .B0(n293), .Y(n288) );
XOR2X1 U317 ( .A(n295), .B(keyIn[4]), .Y(n294) );
OAI21X1 U318 ( .A0(G1036), .A1(n296), .B0(n297), .Y(n295) );
AOI21X1 U319 ( .A0(n298), .A1(n299), .B0(n300), .Y(n287) );
AOI21X1 U320 ( .A0(G132), .A1(G133), .B0(n301), .Y(n300) );
NAND2X1 U321 ( .A(G8), .B(n302), .Y(n299z) );
OAI21X1 U322 ( .A0(G1026), .A1(n303), .B0(n304), .Y(n302) );
OAI21X1 U323 ( .A0(n305), .A1(n306), .B0(n307), .Y(n304) );
AOI21X1 U324 ( .A0(G1026), .A1(n308), .B0(G1021), .Y(n307) );
INVX1 U325 ( .A(n309), .Y(n308) );
AOI21X1 U326 ( .A0(n305), .A1(n306), .B0(n309), .Y(n303) );
AOI21X1 U327 ( .A0(n310), .A1(n309), .B0(n311), .Y(n298) );
AOI21X1 U328 ( .A0(G1033), .A1(G1030), .B0(n312), .Y(n311) );
AOI22X1 U329 ( .A0(n313), .A1(n314), .B0(n315), .B1(n283), .Y(n309) );
AND2X1 U330 ( .A(n306), .B(n305), .Y(n310) );
AOI22X1 U331 ( .A0(n313), .A1(n316), .B0(n315), .B1(n317), .Y(n305z) );
INVX1 U332 ( .A(n312), .Y(n315) );
NAND2X1 U333 ( .A(n318), .B(G8), .Y(n312) );
INVX1 U334 ( .A(n301), .Y(n313) );
NAND2X1 U335 ( .A(G8), .B(n319), .Y(n301) );
AOI21X1 U336 ( .A0(n320), .A1(G1017), .B0(n321), .Y(n306) );
AOI21X1 U337 ( .A0(G2562), .A1(n322), .B0(n323), .Y(n321) );
MX2X1 U338 ( .A(G129), .B(G140), .S0(n318), .Y(n323) );
INVX1 U339 ( .A(n319), .Y(n318) );
INVX1 U340 ( .A(n322), .Y(n320) );
AOI21X1 U341 ( .A0(n324), .A1(n325), .B0(n326), .Y(n322) );
AOI21X1 U342 ( .A0(n327), .A1(n328), .B0(n329), .Y(n326) );
NAND3X1 U343 ( .A(n328), .B(n329), .C(n327), .Y(n325) );
NAND2X1 U344 ( .A(n330), .B(n331), .Y(n327) );
OAI21X1 U345 ( .A0(n331), .A1(n330), .B0(n332), .Y(n328) );
MX2X1 U346 ( .A(n291), .B(n333), .S0(n319), .Y(n332) );
NOR2X1 U347 ( .A(n334), .B(n335), .Y(n330) );
MX2X1 U348 ( .A(G136), .B(G125), .S0(n319), .Y(n334) );
INVX1 U349 ( .A(n336), .Y(n324) );
MX2X1 U350 ( .A(G139), .B(G128), .S0(n319), .Y(n336) );
NAND4X1 U351 ( .A(G30), .B(G2557), .C(n337), .D(n338), .Y(n319) );
AOI22X1 U352 ( .A0(n339), .A1(G138), .B0(G136), .B1(n340), .Y(n285) );
INVX1 U353 ( .A(n290), .Y(n339) );
AOI21X1 U354 ( .A0(n341), .A1(n342), .B0(n293), .Y(n284) );
NAND2X1 U355 ( .A(n343), .B(G30), .Y(n293) );
AOI21X1 U356 ( .A0(n337), .A1(n338), .B0(n344), .Y(n343) );
INVX1 U357 ( .A(G127), .Y(n338) );
OR2X1 U358 ( .A(n340), .B(G136), .Y(n342z) );
AOI22X1 U359 ( .A0(n345), .A1(n297), .B0(n346), .B1(n347), .Y(n341) );
NAND2X1 U360 ( .A(G135), .B(n348), .Y(n297) );
AND2X1 U361 ( .A(n296), .B(G1036), .Y(n345) );
NAND2X1 U362 ( .A(n349), .B(n350), .Y(G2590) );
XOR2X1 U363 ( .A(n351), .B(n352), .Y(n349) );
XOR2X1 U364 ( .A(G1021), .B(G1017), .Y(n352) );
MX2X1 U365 ( .A(n353), .B(n354), .S0(G123), .Y(G2589) );
XOR2X1 U366 ( .A(n355), .B(n351), .Y(n354) );
XOR2X1 U367 ( .A(n356), .B(n357), .Y(n351) );
XOR2X1 U368 ( .A(n358), .B(n359), .Y(n357) );
XOR2X1 U369 ( .A(G1014), .B(n360), .Y(n359) );
XOR2X1 U370 ( .A(n335), .B(n353), .Y(n358) );
XOR2X1 U371 ( .A(n361), .B(n362), .Y(n356) );
XOR2X1 U372 ( .A(G1036), .B(G1033), .Y(n362) );
XOR2X1 U373 ( .A(G1026), .B(G1030), .Y(n361) );
INVX1 U374 ( .A(n363), .Y(n355) );
NAND2X1 U375 ( .A(n364), .B(n350), .Y(G2587) );
INVX1 U376 ( .A(G29), .Y(n350) );
XOR2X1 U377 ( .A(n365), .B(n366), .Y(n364) );
XOR2X1 U378 ( .A(n367), .B(n368), .Y(n366) );
XOR2X1 U379 ( .A(n369), .B(n370), .Y(n368) );
XOR2X1 U380 ( .A(n290), .B(n371), .Y(n370) );
NAND2X1 U381 ( .A(n372), .B(n373), .Y(n371) );
AOI22X1 U382 ( .A0(G84), .A1(n374), .B0(G94), .B1(n375), .Y(n373) );
AOI22X1 U383 ( .A0(G114), .A1(n376), .B0(G104), .B1(n377), .Y(n372) );
XOR2X1 U384 ( .A(n340), .B(n378), .Y(n369) );
XOR2X1 U385 ( .A(n379), .B(n380), .Y(n367) );
XOR2X1 U386 ( .A(n344), .B(n337), .Y(n380) );
XOR2X1 U387 ( .A(G2558), .B(n346), .Y(n379) );
INVX1 U388 ( .A(n348), .Y(n346) );
XOR2X1 U389 ( .A(n353), .B(n381), .Y(G2586) );
NOR2X1 U390 ( .A(G122), .B(n382), .Y(n381) );
XOR2X1 U391 ( .A(n383), .B(n384), .Y(n382) );
NOR2X1 U392 ( .A(n363), .B(n360), .Y(n384) );
NAND2X1 U393 ( .A(n385), .B(n386), .Y(n353) );
AOI22X1 U394 ( .A0(G73), .A1(n387), .B0(G62), .B1(n388), .Y(n386) );
AOI22X1 U395 ( .A0(G41), .A1(n389), .B0(G51), .B1(n390), .Y(n385) );
NAND3X1 U396 ( .A(n391), .B(G9), .C(n392), .Y(G2585) );
MX2X1 U397 ( .A(n393), .B(n394), .S0(G12), .Y(n392) );
NOR2X1 U398 ( .A(n395), .B(n396), .Y(n394) );
NAND4X1 U399 ( .A(n397), .B(n398), .C(n399), .D(n400), .Y(n396) );
XOR2X1 U400 ( .A(n314), .B(G16), .Y(n400) );
XOR2X1 U401 ( .A(n401), .B(G17), .Y(n399) );
XOR2X1 U402 ( .A(n402), .B(G6), .Y(n398) );
XOR2X1 U403 ( .A(n296), .B(G18), .Y(n397) );
NAND4X1 U404 ( .A(n403), .B(n404), .C(n405), .D(n406), .Y(n395) );
XOR2X1 U405 ( .A(n333), .B(G4), .Y(n406) );
NOR2X1 U406 ( .A(n407), .B(n408), .Y(n405) );
XOR2X1 U407 ( .A(G13), .B(G125), .Y(n408) );
XOR2X1 U408 ( .A(G14), .B(G128), .Y(n407) );
XOR2X1 U409 ( .A(n409), .B(G5), .Y(n404) );
XOR2X1 U410 ( .A(n316), .B(G15), .Y(n403) );
NOR2X1 U411 ( .A(n410), .B(n411), .Y(n393) );
NAND4X1 U412 ( .A(n412), .B(n413), .C(n414), .D(n415), .Y(n411) );
XOR2X1 U413 ( .A(n314), .B(G1026), .Y(n415) );
INVX1 U414 ( .A(G131), .Y(n314) );
XOR2X1 U415 ( .A(n401), .B(G1030), .Y(n414) );
INVX1 U416 ( .A(G132), .Y(n401) );
XOR2X1 U417 ( .A(n402), .B(G1033), .Y(n413) );
INVX1 U418 ( .A(G133), .Y(n402) );
XOR2X1 U419 ( .A(n296), .B(G1036), .Y(n412) );
INVX1 U420 ( .A(G134), .Y(n296) );
NAND4X1 U421 ( .A(n416), .B(n417), .C(n418), .D(n419), .Y(n410) );
NOR2X1 U422 ( .A(n420), .B(n421), .Y(n419) );
XOR2X1 U423 ( .A(G1021), .B(G130), .Y(n421) );
XOR2X1 U424 ( .A(G2562), .B(n409), .Y(n420) );
INVX1 U425 ( .A(G129), .Y(n409) );
XOR2X1 U426 ( .A(G125), .B(n383), .Y(n418) );
XOR2X1 U427 ( .A(G128), .B(n329), .Y(n417) );
INVX1 U428 ( .A(G1014), .Y(n329) );
XOR2X1 U429 ( .A(n333), .B(n360), .Y(n416) );
INVX1 U430 ( .A(G126), .Y(n333) );
MX2X1 U431 ( .A(n422), .B(n423), .S0(G23), .Y(n391) );
NOR2X1 U432 ( .A(n424), .B(n425), .Y(n423) );
NAND4X1 U433 ( .A(n426), .B(n427), .C(n428), .D(n429), .Y(n425) );
XOR2X1 U434 ( .A(n291), .B(G20), .Y(n429) );
XOR2X1 U435 ( .A(n430), .B(G21), .Y(n428) );
XOR2X1 U436 ( .A(n317), .B(G26), .Y(n427) );
INVX1 U437 ( .A(G141), .Y(n317) );
XOR2X1 U438 ( .A(n283), .B(G27), .Y(n426) );
INVX1 U439 ( .A(G142), .Y(n283) );
NAND4X1 U440 ( .A(n431), .B(n432), .C(n433), .D(G22), .Y(n424) );
XOR2X1 U441 ( .A(n434), .B(n435), .Y(n433) );
XOR2X1 U442 ( .A(keyIn[3]), .B(G25), .Y(n435) );
XOR2X1 U443 ( .A(n347), .B(G19), .Y(n432) );
XOR2X1 U444 ( .A(n436), .B(G24), .Y(n431) );
NOR2X1 U445 ( .A(n437), .B(n438), .Y(n422) );
NAND4X1 U446 ( .A(n439), .B(n440), .C(n441), .D(n442), .Y(n438) );
XOR2X1 U447 ( .A(n291), .B(n290), .Y(n442) );
NAND2X1 U448 ( .A(n443), .B(n444), .Y(n290) );
AOI22X1 U449 ( .A0(G82), .A1(n374), .B0(G92), .B1(n375), .Y(n444) );
AOI22X1 U450 ( .A0(G112), .A1(n376), .B0(G102), .B1(n377), .Y(n443) );
INVX1 U451 ( .A(G138), .Y(n291) );
XOR2X1 U452 ( .A(n430), .B(n337), .Y(n441) );
INVX1 U453 ( .A(G140), .Y(n430) );
XOR2X1 U454 ( .A(G142), .B(G2558), .Y(n440) );
XOR2X1 U455 ( .A(n344), .B(n445), .Y(n439) );
XOR2X1 U456 ( .A(keyIn[2]), .B(G141), .Y(n445) );
NAND4X1 U457 ( .A(n446), .B(n447), .C(n448), .D(n365), .Y(n437) );
XOR2X1 U458 ( .A(n340), .B(n449), .Y(n448) );
XOR2X1 U459 ( .A(n436), .B(keyIn[1]), .Y(n449) );
INVX1 U460 ( .A(G136), .Y(n436) );
NAND2X1 U461 ( .A(n450), .B(n451), .Y(n340) );
AOI22X1 U462 ( .A0(G83), .A1(n374), .B0(G93), .B1(n375), .Y(n451) );
AOI22X1 U463 ( .A0(G113), .A1(n376), .B0(G103), .B1(n377), .Y(n450) );
XOR2X1 U464 ( .A(n434), .B(n378), .Y(n447) );
NAND2X1 U465 ( .A(n452), .B(n453), .Y(n378z) );
AOI22X1 U466 ( .A0(G81), .A1(n374), .B0(G91), .B1(n375), .Y(n453) );
AOI22X1 U467 ( .A0(G111), .A1(n376), .B0(G101), .B1(n377), .Y(n452) );
INVX1 U468 ( .A(G139), .Y(n434) );
XOR2X1 U469 ( .A(n347), .B(n348), .Y(n446) );
NAND2X1 U470 ( .A(n454), .B(n455), .Y(n348) );
AOI22X1 U471 ( .A0(G75), .A1(n374), .B0(G85), .B1(n375), .Y(n455) );
AOI22X1 U472 ( .A0(G105), .A1(n376), .B0(G95), .B1(n377), .Y(n454) );
INVX1 U473 ( .A(G135), .Y(n347) );
XOR2X1 U474 ( .A(n456), .B(n457), .Y(G2583) );
XOR2X1 U475 ( .A(n458), .B(n459), .Y(n457) );
XOR2X1 U476 ( .A(n460), .B(n461), .Y(n459) );
XOR2X1 U477 ( .A(G129), .B(G128), .Y(n461) );
XOR2X1 U478 ( .A(G132), .B(G131), .Y(n460) );
XOR2X1 U479 ( .A(n462), .B(n463), .Y(n458) );
XOR2X1 U480 ( .A(G135), .B(G133), .Y(n463) );
XOR2X1 U481 ( .A(G156), .B(G136), .Y(n462) );
XOR2X1 U482 ( .A(n316), .B(G134), .Y(n456) );
INVX1 U483 ( .A(G130), .Y(n316) );
NAND2X1 U484 ( .A(G10), .B(n464), .Y(G2581) );
XOR2X1 U485 ( .A(n465), .B(n466), .Y(n464) );
XOR2X1 U486 ( .A(G152), .B(n467), .Y(n466) );
XOR2X1 U487 ( .A(n468), .B(n469), .Y(n467) );
XOR2X1 U488 ( .A(n470), .B(n471), .Y(n469) );
XOR2X1 U489 ( .A(G126), .B(G125), .Y(n471) );
XOR2X1 U490 ( .A(G149), .B(G148), .Y(n470) );
XOR2X1 U491 ( .A(n472), .B(n473), .Y(n468) );
XOR2X1 U492 ( .A(G151), .B(G150), .Y(n473) );
XOR2X1 U493 ( .A(G155), .B(G154), .Y(n472) );
XOR2X1 U494 ( .A(keyIn[0]), .B(G153), .Y(n465) );
NAND2X1 U495 ( .A(n474), .B(n475), .Y(G2580) );
INVX1 U496 ( .A(G144), .Y(n475) );
XOR2X1 U497 ( .A(n365), .B(G143), .Y(n474) );
NAND2X1 U498 ( .A(n476), .B(n477), .Y(n365) );
AOI22X1 U499 ( .A0(G77), .A1(n374), .B0(G87), .B1(n375), .Y(n477) );
AOI22X1 U500 ( .A0(G107), .A1(n376), .B0(G97), .B1(n377), .Y(n476) );
MX2X1 U501 ( .A(n383), .B(n363), .S0(G123), .Y(G2579) );
OAI21X1 U502 ( .A0(G122), .A1(n363), .B0(n331), .Y(G2577) );
NOR2X1 U503 ( .A(G118), .B(n360), .Y(n363) );
MX2X1 U504 ( .A(G1014), .B(G2561), .S0(G123), .Y(G2576) );
MX2X1 U505 ( .A(n331), .B(G1017), .S0(G123), .Y(G2574) );
INVX1 U506 ( .A(n360), .Y(n331) );
NAND2X1 U507 ( .A(n478), .B(n479), .Y(n360) );
AOI22X1 U508 ( .A0(G72), .A1(n387), .B0(G61), .B1(n388), .Y(n479) );
AOI22X1 U509 ( .A0(G40), .A1(n389), .B0(G50), .B1(n390), .Y(n478) );
INVX1 U510 ( .A(n480), .Y(G2565) );
AOI21X1 U511 ( .A0(G3), .A1(G1), .B0(n481), .Y(n480) );
NAND2X1 U512 ( .A(G28), .B(n482), .Y(G2564) );
INVX1 U513 ( .A(n481), .Y(n482) );
NAND3X1 U514 ( .A(n273), .B(n483), .C(G116), .Y(n481) );
INVX1 U515 ( .A(G121), .Y(n483) );
NAND2X1 U516 ( .A(G122), .B(n383), .Y(G2563) );
INVX1 U517 ( .A(n335), .Y(n383) );
NAND2X1 U518 ( .A(n484), .B(n485), .Y(n335) );
AOI22X1 U519 ( .A0(G63), .A1(n387), .B0(G52), .B1(n388), .Y(n485) );
AOI22X1 U520 ( .A0(G31), .A1(n389), .B0(G42), .B1(n390), .Y(n484) );
INVX1 U521 ( .A(G1017), .Y(G2562) );
INVX1 U522 ( .A(G1021), .Y(G2561) );
INVX1 U523 ( .A(G1026), .Y(G2560) );
INVX1 U524 ( .A(n337), .Y(G2559) );
NAND2X1 U525 ( .A(n486), .B(n487), .Y(n337) );
AOI22X1 U526 ( .A0(G80), .A1(n374), .B0(G90), .B1(n375), .Y(n487) );
AOI22X1 U527 ( .A0(G110), .A1(n376), .B0(G100), .B1(n377), .Y(n486) );
AND2X1 U528 ( .A(n488), .B(n489), .Y(G2558) );
AOI22X1 U529 ( .A0(G78), .A1(n374), .B0(G88), .B1(n375), .Y(n489) );
AOI22X1 U530 ( .A0(G108), .A1(n376), .B0(G98), .B1(n377), .Y(n488) );
INVX1 U531 ( .A(n344), .Y(G2557) );
NAND2X1 U532 ( .A(n490), .B(n491), .Y(n344) );
AOI22X1 U533 ( .A0(G79), .A1(n374), .B0(G89), .B1(n375), .Y(n491) );
NOR2X1 U534 ( .A(G145), .B(G146), .Y(n375) );
NOR2X1 U535 ( .A(n492), .B(G145), .Y(n374) );
AOI22X1 U536 ( .A0(G109), .A1(n376), .B0(G99), .B1(n377), .Y(n490z) );
NOR2X1 U537 ( .A(n493), .B(G146), .Y(n377) );
NOR2X1 U538 ( .A(n493), .B(n492), .Y(n376) );
INVX1 U539 ( .A(G146), .Y(n492) );
INVX1 U540 ( .A(G145), .Y(n493) );
INVX1 U541 ( .A(n273), .Y(G2556) );
AOI22X1 U542 ( .A0(G147), .A1(n494), .B0(G119), .B1(n495), .Y(n273) );
OR2X1 U543 ( .A(n495), .B(n494), .Y(G2555) );
NAND4X1 U544 ( .A(G32), .B(G106), .C(G64), .D(G76), .Y(n494) );
NAND4X1 U545 ( .A(G43), .B(G53), .C(G96), .D(G86), .Y(n495) );
NAND2X1 U546 ( .A(G147), .B(n496), .Y(G2553) );
NAND2X1 U547 ( .A(G119), .B(n496), .Y(G2552) );
INVX1 U548 ( .A(G2551), .Y(n496) );
NAND2X1 U549 ( .A(G7), .B(G121), .Y(G2551) );
AND2X1 U550 ( .A(G74), .B(G2531), .Y(G2550) );
NAND3X1 U551 ( .A(G11), .B(G121), .C(G2), .Y(G2548) );
NAND4X1 U552 ( .A(G139), .B(G140), .C(G141), .D(G142), .Y(G2547) );
INVX1 U553 ( .A(G86), .Y(G2546) );
XOR2X1 U554 ( .A(keyIn[7]), .B(G43), .Y(G2545) );
INVX1 U555 ( .A(G96), .Y(G2544) );
INVX1 U556 ( .A(G53), .Y(G2543) );
INVX1 U557 ( .A(G76), .Y(G2542) );
INVX1 U558 ( .A(G64), .Y(G2541) );
INVX1 U559 ( .A(G106), .Y(G2540) );
INVX1 U560 ( .A(G32), .Y(G2539) );
XOR2X1 U561 ( .A(keyIn[5]), .B(G137), .Y(G2538) );
INVX1 U562 ( .A(G124), .Y(G2534) );
INVX1 U563 ( .A(G115), .Y(G2531) );
NAND2X1 U564 ( .A(n497), .B(n498), .Y(G1036) );
AOI22X1 U565 ( .A0(G65), .A1(n387), .B0(G54), .B1(n388), .Y(n498) );
AOI22X1 U566 ( .A0(G33), .A1(n389), .B0(G44), .B1(n390), .Y(n497) );
NAND2X1 U567 ( .A(n499), .B(n500), .Y(G1033) );
AOI22X1 U568 ( .A0(G66), .A1(n387), .B0(G55), .B1(n388), .Y(n500) );
AOI22X1 U569 ( .A0(G34), .A1(n389), .B0(G45), .B1(n390), .Y(n499) );
NAND2X1 U570 ( .A(n501), .B(n502), .Y(G1030) );
AOI21X1 U571 ( .A0(G35), .A1(n389), .B0(n390), .Y(n502) );
AOI22X1 U572 ( .A0(G67), .A1(G117), .B0(G56), .B1(n503), .Y(n501) );
NAND2X1 U573 ( .A(n504), .B(n505), .Y(G1026) );
AOI22X1 U574 ( .A0(G68), .A1(n387), .B0(G57), .B1(n388), .Y(n505) );
AOI22X1 U575 ( .A0(G36), .A1(n389), .B0(G46), .B1(n390), .Y(n504) );
NAND2X1 U576 ( .A(n506), .B(n507), .Y(G1021) );
AOI22X1 U577 ( .A0(G69), .A1(n387), .B0(G58), .B1(n388), .Y(n507) );
AOI22X1 U578 ( .A0(G37), .A1(n389), .B0(G47), .B1(n390), .Y(n506) );
NAND2X1 U579 ( .A(n508), .B(n509), .Y(G1017z) );
AOI22X1 U580 ( .A0(G70), .A1(n387), .B0(G59), .B1(n388), .Y(n509) );
AOI22X1 U581 ( .A0(G38), .A1(n389), .B0(G48), .B1(n390), .Y(n508) );
NAND2X1 U582 ( .A(n510), .B(n511), .Y(G1014) );
XOR2X1 U583 ( .A(keyIn[6]), .B(n512), .Y(n511) );
AOI22X1 U584 ( .A0(G60), .A1(n388), .B0(G71), .B1(n387), .Y(n512) );
NOR2X1 U585 ( .A(n503), .B(n513), .Y(n387) );
NOR2X1 U586 ( .A(G117), .B(G120), .Y(n388) );
AOI22X1 U587 ( .A0(G39), .A1(n389), .B0(G49), .B1(n390), .Y(n510) );
NOR2X1 U588 ( .A(n513), .B(G120), .Y(n390) );
INVX1 U589 ( .A(G117), .Y(n513) );
NOR2X1 U590 ( .A(n503), .B(G117), .Y(n389) );
INVX1 U591 ( .A(G120), .Y(n503) );
  XOR2X1 enc2XOR2X10 ( .A(keyInPseudo[5]), .B(G2533z), .Y(G2533) );
  XOR2X1 enc2XOR2X11 ( .A(keyInPseudo[3]), .B(n305z), .Y(n305) );
  XOR2X1 enc2XOR2X12 ( .A(keyInPseudo[7]), .B(G1017z), .Y(G1017) );
  XOR2X1 enc2XOR2X13 ( .A(keyInPseudo[6]), .B(G2569z), .Y(G2569z_inv_wire) );
  INVX1 inv0inv( .A(G2569z_inv_wire), .Y(G2569) );
  XOR2X1 enc2XOR2X14 ( .A(keyInPseudo[1]), .B(n299z), .Y(n299) );
  XOR2X1 enc2XOR2X15 ( .A(keyInPseudo[4]), .B(n342z), .Y(n342) );
  XOR2X1 enc2XOR2X16 ( .A(keyInPseudo[2]), .B(n490z), .Y(n490) );
  XOR2X1 enc2XOR2X17 ( .A(keyInPseudo[0]), .B(n378z), .Y(n378z_inv_wire) );
  INVX1 inv1inv( .A(n378z_inv_wire), .Y(n378) );
endmodule